module inverseAdd_Round_Key(
  input  [127:0] in,
  input  [127:0] key,
  output [127:0] out
  );
  //same implementation of add round key
Add_Round_Key inverse(in,key,out);
endmodule
