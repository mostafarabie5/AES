module inverse_ShiftRows_tb();

reg [0:127] in;
wire [0:127] out;	


inverse_ShiftRows m (in,out);


initial begin
	$monitor("input= %H , output= %h",in,out);
	in = 128'h_d4bf5d30_e0b452ae_b84111f1_1e2798e5;
	#10;
	in = 128'h_49db873b_45395389_7f02d2f1_77de961a;
	#10;
	in = 128'h_acc1d6b8_efb55a7b_1323cfdf_457311b5;
end
endmodule
